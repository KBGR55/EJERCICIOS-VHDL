----------------------------------------------------------------------------------
-- Karen Brigith Gonzaga Rivas
-- Create Date:    18:54:40 05/23/2022 
-- Pregunta : 1.9
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity and_gate is
    Port ( A,B : in  STD_LOGIC;
           C : out  STD_LOGIC);
end and_gate;

architecture Behavioral of and_gate is

begin


end Behavioral;

