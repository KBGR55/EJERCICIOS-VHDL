----------------------------------------------------------------------------------
-- Create Date:    19:25:38 05/23/2022 
-- Karen Brigith Gonzaga Rivas
-- Pregunta : 1.11
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Promedio_01 is
    Port ( A,B : in  STD_LOGIC_VECTOR (2 downto 0);
           C : out  STD_LOGIC_VECTOR (2 downto 0));
end Promedio_01;

architecture Behavioral of Promedio_01 is

begin

end Behavioral;