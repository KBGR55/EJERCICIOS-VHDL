----------------------------------------------------------------------------------
-- Create Date:    21:55:16 05/23/2022 
-- Karen Brigith Gonzaga Rivas
-- Pregunta : 1.16
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX_VECTOR4_1 is
    Port ( E0,E1,E2,E3 : in  STD_LOGIC_VECTOR (3 downto 0);
           S0,S1 : in  STD_LOGIC_VECTOR (3 downto 0);
           F : out  STD_LOGIC);
end MUX_VECTOR4_1;

architecture Behavioral of MUX_VECTOR4_1 is

begin

end Behavioral;