----------------------------------------------------------------------------------
-- Create Date:    21:52:17 05/23/2022 
-- Karen Brigith Gonzaga Rivas
-- Pregunta : 1.15
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX4_1 is
    Port ( E0,E1,E2,E3 : in  STD_LOGIC;
           S0,S1 : in  STD_LOGIC;
           F : out  STD_LOGIC);
end MUX4_1;

architecture Behavioral of MUX4_1 is

begin

end Behavioral;