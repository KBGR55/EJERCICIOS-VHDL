----------------------------------------------------------------------------------
-- Create Date:    19:27:57 05/23/2022 
-- Karen Brigith Gonzaga Rivas
-- Pregunta : 1.11
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Promedio_02 is
    Port ( A,B : in  STD_LOGIC_VECTOR (0 to 3);
           C : out  STD_LOGIC_VECTOR (0 to 3));
end Promedio_02;

architecture Behavioral of Promedio_02 is

begin

end Behavioral;