----------------------------------------------------------------------------------
-- Karen Gonzaga Rivas
-- Create Date:    18:54:40 05/23/2022 
-- Pregunta : 1.8 
---------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ejemplo is
    Port ( X1,X2 : in  STD_LOGIC;
           fa,fb : out  STD_LOGIC);
end ejemplo;

architecture Behavioral of ejemplo is

begin

end Behavioral;