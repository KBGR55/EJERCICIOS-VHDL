----------------------------------------------------------------------------------
-- Karen Brigith Gonzaga Rivas
-- Create Date:    18:59:38 05/23/2022 
-- Pregunta : 1.9
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Proyecto is
    Port ( P0,P1,P2 : in  STD_LOGIC;
			  X : buffer STD_LOGIC;
           A0,A1 : out  STD_LOGIC);
end Proyecto;

architecture Behavioral of Proyecto is

begin

end Behavioral;